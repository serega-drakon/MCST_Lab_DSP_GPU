module Control (

);



endmodule
module ALU (

);



endmodule : ALU
module GPU(
    input wire clk,
    input wire reset
);



endmodule
module Core #()(
    input wire init_R0_flag

    );



endmodule
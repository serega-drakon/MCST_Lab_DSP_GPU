`ifndef CONSTANTS
`define CONSTANTS

`define INSN_COUNT 16
`define INSN_SIZE 2
`define INSN_PTR_SIZE 4
`define INSN_OPC_SIZE 4
`define REG_COUNT 16
`define REG_PTR_SIZE 4
`define REG_SIZE 8
`define CORE_ID_SIZE 4
`define ADDR_SIZE (`CORE_ID_SIZE + `REG_SIZE) //ну по смыслу близко)

`endif //CONSTANTS
module RegisterFile (

);
    localparam REG_SIZE = `REG_SIZE;
    localparam REG_PTR_SIZE = `REG_PTR_SIZE;


endmodule
`define INSN_COUNT 16
`define INSN_SIZE 2
`define INSN_PTR_SIZE 4
`define REG_COUNT 16
`define REG_PTR_SIZE 4
`define REG_SIZE 8
`define ADDR_SIZE 12

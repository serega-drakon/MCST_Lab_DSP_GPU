`include "Inc/Instruction Set.vh"
`include "Inc/Constants.vh"

module ALU (

);



endmodule : ALU